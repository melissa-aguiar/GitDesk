library verilog;
use verilog.vl_types.all;
entity proc_fix_tb is
end proc_fix_tb;
