library verilog;
use verilog.vl_types.all;
entity proc_v1_tb is
end proc_v1_tb;
