library verilog;
use verilog.vl_types.all;
entity proc_float_tb is
end proc_float_tb;
