module multicore_tb();

reg         		 clk;//, rst;
wire			[ 1:0] req_in0, req_in1;//, req_in2, req_in3, req_in4, req_in5, req_in6, req_in7, req_in8, req_in9, req_in10, req_in11, req_in12, req_in13, req_in14, req_in15, req_in16, req_in17, req_in18, req_in19, req_in20, req_in21, req_in22, req_in23, req_in24, req_in25, req_in26, req_in27, req_in28, req_in29, req_in30, req_in31, req_in32, req_in33, req_in34, req_in35, req_in36, req_in37, req_in38, req_in39, req_in40, req_in41, req_in42, req_in43, req_in44, req_in45, req_in46, req_in47, req_in48, req_in49, req_in50, req_in51, req_in52, req_in53, req_in54, req_in55, req_in56, req_in57, req_in58, req_in59, req_in60, req_in61, req_in62, req_in63, req_in64, req_in65, req_in66, req_in67, req_in68, req_in69, req_in70, req_in71, req_in72, req_in73, req_in74, req_in75, req_in76, req_in77, req_in78, req_in79, req_in80, req_in81, req_in82, req_in83, req_in84, req_in85, req_in86, req_in87, req_in88, req_in89, req_in90, req_in91, req_in92, req_in93, req_in94, req_in95, req_in96, req_in97, req_in98, req_in99, req_in100, req_in101, req_in102, req_in103, req_in104, req_in105, req_in106, req_in107, req_in108, req_in109, req_in110, req_in111, req_in112, req_in113, req_in114, req_in115, req_in116, req_in117, req_in118, req_in119, req_in120, req_in121, req_in122, req_in123, req_in124, req_in125, req_in126, req_in127, req_in128, req_in129, req_in130, req_in131, req_in132, req_in133, req_in134, req_in135, req_in136, req_in137, req_in138, req_in139;
reg signed  [28:0] in;
wire signed [28:0] io_out0, io_out1;//, io_out2, io_out3, io_out4, io_out5, io_out6, io_out7, io_out8, io_out9, io_out10, io_out11, io_out12, io_out13, io_out14, io_out15, io_out16, io_out17, io_out18, io_out19, io_out20, io_out21, io_out22, io_out23, io_out24, io_out25, io_out26, io_out27, io_out28, io_out29, io_out30, io_out31, io_out32, io_out33, io_out34, io_out35, io_out36, io_out37, io_out38, io_out39, io_out40, io_out41, io_out42, io_out43, io_out44, io_out45, io_out46, io_out47, io_out48, io_out49, io_out50, io_out51, io_out52, io_out53, io_out54, io_out55, io_out56, io_out57, io_out58, io_out59, io_out60, io_out61, io_out62, io_out63, io_out64, io_out65, io_out66, io_out67, io_out68, io_out69, io_out70, io_out71, io_out72, io_out73, io_out74, io_out75, io_out76, io_out77, io_out78, io_out79, io_out80, io_out81, io_out82, io_out83, io_out84, io_out85, io_out86, io_out87, io_out88, io_out89, io_out90, io_out91, io_out92, io_out93, io_out94, io_out95, io_out96, io_out97, io_out98, io_out99, io_out100, io_out101, io_out102, io_out103, io_out104, io_out105, io_out106, io_out107, io_out108, io_out109, io_out110, io_out111, io_out112, io_out113, io_out114, io_out115, io_out116, io_out117, io_out118, io_out119, io_out120, io_out121, io_out122, io_out123, io_out124, io_out125, io_out126, io_out127, io_out128, io_out129, io_out130, io_out131, io_out132, io_out133, io_out134, io_out135, io_out136, io_out137, io_out138, io_out139;
wire 			[ 1:0] out_en0, out_en1;//, out_en2, out_en3, out_en4, out_en5, out_en6, out_en7, out_en8, out_en9, out_en10, out_en11, out_en12, out_en13, out_en14, out_en15, out_en16, out_en17, out_en18, out_en19, out_en20, out_en21, out_en22, out_en23, out_en24, out_en25, out_en26, out_en27, out_en28, out_en29, out_en30, out_en31, out_en32, out_en33, out_en34, out_en35, out_en36, out_en37, out_en38, out_en39, out_en40, out_en41, out_en42, out_en43, out_en44, out_en45, out_en46, out_en47, out_en48, out_en49, out_en50, out_en51, out_en52, out_en53, out_en54, out_en55, out_en56, out_en57, out_en58, out_en59, out_en60, out_en61, out_en62, out_en63, out_en64, out_en65, out_en66, out_en67, out_en68, out_en69, out_en70, out_en71, out_en72, out_en73, out_en74, out_en75, out_en76, out_en77, out_en78, out_en79, out_en80, out_en81, out_en82, out_en83, out_en84, out_en85, out_en86, out_en87, out_en88, out_en89, out_en90, out_en91, out_en92, out_en93, out_en94, out_en95, out_en96, out_en97, out_en98, out_en99, out_en100, out_en101, out_en102, out_en103, out_en104, out_en105, out_en106, out_en107, out_en108, out_en109, out_en110, out_en111, out_en112, out_en113, out_en114, out_en115, out_en116, out_en117, out_en118, out_en119, out_en120, out_en121, out_en122, out_en123, out_en124, out_en125, out_en126, out_en127, out_en128, out_en129, out_en130, out_en131, out_en132, out_en133, out_en134, out_en135, out_en136, out_en137, out_en138, out_en139;
integer 				 data_file, scan_file, my_output;



initial begin 
	//data_file = $fopen("signalN_48b7e_30.txt", "r");
	data_file = $fopen("signalN.txt", "r");
	my_output = $fopen("myoutput.txt", "w");
	scan_file = $fscanf(data_file, "%d\n", in);
	clk = 0;
	//rst  = 1;
	//#1 rst = 0;
end

always #1000 clk = ~clk;



always @(posedge clk) begin
	if ((req_in0 || req_in1) == 1'd1) //|| req_in2 || req_in3 || req_in4 || req_in5 || req_in6 || req_in7 || req_in8 || req_in9 || req_in10 || req_in11 || req_in12 || req_in13 || req_in14 || req_in15 || req_in16 || req_in17 || req_in18 || req_in19 || req_in20 || req_in21 || req_in22 || req_in23 || req_in24 || req_in25 || req_in26 || req_in27 || req_in28 || req_in29 || req_in30 || req_in31 || req_in32 || req_in33 || req_in34 || req_in35 || req_in36 || req_in37 || req_in38 || req_in39 || req_in40 || req_in41 || req_in42 || req_in43 || req_in44 || req_in45 || req_in46 || req_in47 || req_in48 || req_in49 || req_in50 || req_in51 || req_in52 || req_in53 || req_in54 || req_in55 || req_in56 || req_in57 || req_in58 || req_in59 || req_in60 || req_in61 || req_in62 || req_in63 || req_in64 || req_in65 || req_in66 || req_in67 || req_in68 || req_in69 || req_in70 || req_in71 || req_in72 || req_in73 || req_in74 || req_in75 || req_in76 || req_in77 || req_in78 || req_in79 || req_in80 || req_in81 || req_in82 || req_in83 || req_in84 || req_in85 || req_in86 || req_in87 || req_in88 || req_in89 || req_in90 || req_in91 || req_in92 || req_in93 || req_in94 || req_in95 || req_in96 || req_in97 || req_in98 || req_in99 || req_in100 || req_in101 || req_in102 || req_in103 || req_in104 || req_in105 || req_in106 || req_in107 || req_in108 || req_in109 || req_in110 || req_in111 || req_in112 || req_in113 || req_in114 || req_in115 || req_in116 || req_in117 || req_in118 || req_in119 || req_in120 || req_in121 || req_in122 || req_in123 || req_in124 || req_in125 || req_in126 || req_in127 || req_in128 || req_in129 || req_in130 || req_in131 || req_in132 || req_in133 || req_in134 || req_in135 || req_in136 || req_in137 || req_in138 || req_in139) == 1'd1)
		scan_file = $fscanf(data_file, "%d\n", in);
end

always @ (posedge clk) begin
	//if ((out_en || out_en0 || out_en1 || out_en2 || out_en3 || out_en4 || out_en5 || out_en6 || out_en7 || out_en8 || out_en9 || out_en10 || out_en11 || out_en12 || out_en13 || out_en14 || out_en15 || out_en16 || out_en17 || out_en18 || out_en19 || out_en20 || out_en21 || out_en22 || out_en23 || out_en24 || out_en25 || out_en26 || out_en27 || out_en28 || out_en29 || out_en30 || out_en31 || out_en32 || out_en33 || out_en34 || out_en35 || out_en36 || out_en37 || out_en38 || out_en39 || out_en40 || out_en41 || out_en42 || out_en43 || out_en44 || out_en45 || out_en46 || out_en47 || out_en48 || out_en49 || out_en50 || out_en51 || out_en52 || out_en53 || out_en54 || out_en55 || out_en56 || out_en57 || out_en58 || out_en59 || out_en60 || out_en61 || out_en62 || out_en63 || out_en64 || out_en65 || out_en66 || out_en67 || out_en68 || out_en69 || out_en70 || out_en71 || out_en72 || out_en73 || out_en74 || out_en75 || out_en76 || out_en77 || out_en78 || out_en79 || out_en80 || out_en81 || out_en82 || out_en83 || out_en84 || out_en85 || out_en86 || out_en87 || out_en88 || out_en89 || out_en90 || out_en91 || out_en92 || out_en93 || out_en94 || out_en95 || out_en96 || out_en97 || out_en98 || out_en99 || out_en100 || out_en101 || out_en102 || out_en103 || out_en104 || out_en105 || out_en106 || out_en107 || out_en108 || out_en109 || out_en110 || out_en111 || out_en112 || out_en113 || out_en114 || out_en115 || out_en116 || out_en117 || out_en118 || out_en119 || out_en120 || out_en121 || out_en122 || out_en123 || out_en124 || out_en125 || out_en126 || out_en127 || out_en128 || out_en129 || out_en130 || out_en131 || out_en132 || out_en133 || out_en134 || out_en135 || out_en136 || out_en137 || out_en138 || out_en139 || out_en140 || out_en141 || out_en142 || out_en143 || out_en144 || out_en145 || out_en146 || out_en147 || out_en148 || out_en149 || out_en150 || out_en151 || out_en152 || out_en153 || out_en154 || out_en155 || out_en156 || out_en157 || out_en158 || out_en159 || out_en160 || out_en161 || out_en162 || out_en163 || out_en164 || out_en165 || out_en166 || out_en167 || out_en168 || out_en169 || out_en170) == 1'd1)
	if (out_en0 == 1'd1) $fwrite(my_output, "%d\n", io_out0);
	if (out_en1 == 1'd1) $fwrite(my_output, "%d\n", io_out1);
	//if (out_en2 == 1'd1) $fwrite(my_output, "%d\n", io_out2);
	//if (out_en3 == 1'd1) $fwrite(my_output, "%d\n", io_out3);
	//if (out_en4 == 1'd1) $fwrite(my_output, "%d\n", io_out4);
	//if (out_en5 == 1'd1) $fwrite(my_output, "%d\n", io_out5);
	//if (out_en6 == 1'd1) $fwrite(my_output, "%d\n", io_out6);
	//if (out_en7 == 1'd1) $fwrite(my_output, "%d\n", io_out7);
	//if (out_en8 == 1'd1) $fwrite(my_output, "%d\n", io_out8);
	//if (out_en9 == 1'd1) $fwrite(my_output, "%d\n", io_out9);
	//if (out_en10 == 1'd1) $fwrite(my_output, "%d\n", io_out10);
	//if (out_en11 == 1'd1) $fwrite(my_output, "%d\n", io_out11);
	//if (out_en12 == 1'd1) $fwrite(my_output, "%d\n", io_out12);
	//if (out_en13 == 1'd1) $fwrite(my_output, "%d\n", io_out13);
	//if (out_en14 == 1'd1) $fwrite(my_output, "%d\n", io_out14);
	//if (out_en15 == 1'd1) $fwrite(my_output, "%d\n", io_out15);
	//if (out_en16 == 1'd1) $fwrite(my_output, "%d\n", io_out16);
	//if (out_en17 == 1'd1) $fwrite(my_output, "%d\n", io_out17);
	//if (out_en18 == 1'd1) $fwrite(my_output, "%d\n", io_out18);
	//if (out_en19 == 1'd1) $fwrite(my_output, "%d\n", io_out19);
	//if (out_en20 == 1'd1) $fwrite(my_output, "%d\n", io_out20);
	//if (out_en21 == 1'd1) $fwrite(my_output, "%d\n", io_out21);
	//if (out_en22 == 1'd1) $fwrite(my_output, "%d\n", io_out22);
	//if (out_en23 == 1'd1) $fwrite(my_output, "%d\n", io_out23);
	//if (out_en24 == 1'd1) $fwrite(my_output, "%d\n", io_out24);
	//if (out_en25 == 1'd1) $fwrite(my_output, "%d\n", io_out25);
	//if (out_en26 == 1'd1) $fwrite(my_output, "%d\n", io_out26);
	//if (out_en27 == 1'd1) $fwrite(my_output, "%d\n", io_out27);
	//if (out_en28 == 1'd1) $fwrite(my_output, "%d\n", io_out28);
	//if (out_en29 == 1'd1) $fwrite(my_output, "%d\n", io_out29);
	//if (out_en30 == 1'd1) $fwrite(my_output, "%d\n", io_out30);
	//if (out_en31 == 1'd1) $fwrite(my_output, "%d\n", io_out31);
	//if (out_en32 == 1'd1) $fwrite(my_output, "%d\n", io_out32);
	//if (out_en33 == 1'd1) $fwrite(my_output, "%d\n", io_out33);
	//if (out_en34 == 1'd1) $fwrite(my_output, "%d\n", io_out34);
	//if (out_en35 == 1'd1) $fwrite(my_output, "%d\n", io_out35);
	//if (out_en36 == 1'd1) $fwrite(my_output, "%d\n", io_out36);
	//if (out_en37 == 1'd1) $fwrite(my_output, "%d\n", io_out37);
	//if (out_en38 == 1'd1) $fwrite(my_output, "%d\n", io_out38);
	//if (out_en39 == 1'd1) $fwrite(my_output, "%d\n", io_out39);
	//if (out_en40 == 1'd1) $fwrite(my_output, "%d\n", io_out40);
	//if (out_en41 == 1'd1) $fwrite(my_output, "%d\n", io_out41);
	//if (out_en42 == 1'd1) $fwrite(my_output, "%d\n", io_out42);
	//if (out_en43 == 1'd1) $fwrite(my_output, "%d\n", io_out43);
	//if (out_en44 == 1'd1) $fwrite(my_output, "%d\n", io_out44);
	//if (out_en45 == 1'd1) $fwrite(my_output, "%d\n", io_out45);
	//if (out_en46 == 1'd1) $fwrite(my_output, "%d\n", io_out46);
	//if (out_en47 == 1'd1) $fwrite(my_output, "%d\n", io_out47);
	//if (out_en48 == 1'd1) $fwrite(my_output, "%d\n", io_out48);
	//if (out_en49 == 1'd1) $fwrite(my_output, "%d\n", io_out49);
	//if (out_en50 == 1'd1) $fwrite(my_output, "%d\n", io_out50);
	//if (out_en51 == 1'd1) $fwrite(my_output, "%d\n", io_out51);
	//if (out_en52 == 1'd1) $fwrite(my_output, "%d\n", io_out52);
	//if (out_en53 == 1'd1) $fwrite(my_output, "%d\n", io_out53);
	//if (out_en54 == 1'd1) $fwrite(my_output, "%d\n", io_out54);
	//if (out_en55 == 1'd1) $fwrite(my_output, "%d\n", io_out55);
	//if (out_en56 == 1'd1) $fwrite(my_output, "%d\n", io_out56);
	//if (out_en57 == 1'd1) $fwrite(my_output, "%d\n", io_out57);
	//if (out_en58 == 1'd1) $fwrite(my_output, "%d\n", io_out58);
	//if (out_en59 == 1'd1) $fwrite(my_output, "%d\n", io_out59);
	//if (out_en60 == 1'd1) $fwrite(my_output, "%d\n", io_out60);
	//if (out_en61 == 1'd1) $fwrite(my_output, "%d\n", io_out61);
	//if (out_en62 == 1'd1) $fwrite(my_output, "%d\n", io_out62);
	//if (out_en63 == 1'd1) $fwrite(my_output, "%d\n", io_out63);
	//if (out_en64 == 1'd1) $fwrite(my_output, "%d\n", io_out64);
	//if (out_en65 == 1'd1) $fwrite(my_output, "%d\n", io_out65);
	//if (out_en66 == 1'd1) $fwrite(my_output, "%d\n", io_out66);
	//if (out_en67 == 1'd1) $fwrite(my_output, "%d\n", io_out67);
	//if (out_en68 == 1'd1) $fwrite(my_output, "%d\n", io_out68);
	//if (out_en69 == 1'd1) $fwrite(my_output, "%d\n", io_out69);
	//if (out_en70 == 1'd1) $fwrite(my_output, "%d\n", io_out70);
	//if (out_en71 == 1'd1) $fwrite(my_output, "%d\n", io_out71);
	//if (out_en72 == 1'd1) $fwrite(my_output, "%d\n", io_out72);
	//if (out_en73 == 1'd1) $fwrite(my_output, "%d\n", io_out73);
	//if (out_en74 == 1'd1) $fwrite(my_output, "%d\n", io_out74);
	//if (out_en75 == 1'd1) $fwrite(my_output, "%d\n", io_out75);
	//if (out_en76 == 1'd1) $fwrite(my_output, "%d\n", io_out76);
	//if (out_en77 == 1'd1) $fwrite(my_output, "%d\n", io_out77);
	//if (out_en78 == 1'd1) $fwrite(my_output, "%d\n", io_out78);
	//if (out_en79 == 1'd1) $fwrite(my_output, "%d\n", io_out79);
	//if (out_en80 == 1'd1) $fwrite(my_output, "%d\n", io_out80);
	//if (out_en81 == 1'd1) $fwrite(my_output, "%d\n", io_out81);
	//if (out_en82 == 1'd1) $fwrite(my_output, "%d\n", io_out82);
	//if (out_en83 == 1'd1) $fwrite(my_output, "%d\n", io_out83);
	//if (out_en84 == 1'd1) $fwrite(my_output, "%d\n", io_out84);
	//if (out_en85 == 1'd1) $fwrite(my_output, "%d\n", io_out85);
	//if (out_en86 == 1'd1) $fwrite(my_output, "%d\n", io_out86);
	//if (out_en87 == 1'd1) $fwrite(my_output, "%d\n", io_out87);
	//if (out_en88 == 1'd1) $fwrite(my_output, "%d\n", io_out88);
	//if (out_en89 == 1'd1) $fwrite(my_output, "%d\n", io_out89);
	//if (out_en90 == 1'd1) $fwrite(my_output, "%d\n", io_out90);
	//if (out_en91 == 1'd1) $fwrite(my_output, "%d\n", io_out91);
	//if (out_en92 == 1'd1) $fwrite(my_output, "%d\n", io_out92);
	//if (out_en93 == 1'd1) $fwrite(my_output, "%d\n", io_out93);
	//if (out_en94 == 1'd1) $fwrite(my_output, "%d\n", io_out94);
	//if (out_en95 == 1'd1) $fwrite(my_output, "%d\n", io_out95);
	//if (out_en96 == 1'd1) $fwrite(my_output, "%d\n", io_out96);
	//if (out_en97 == 1'd1) $fwrite(my_output, "%d\n", io_out97);
	//if (out_en98 == 1'd1) $fwrite(my_output, "%d\n", io_out98);
	//if (out_en99 == 1'd1) $fwrite(my_output, "%d\n", io_out99);
	//if (out_en100 == 1'd1) $fwrite(my_output, "%d\n", io_out100);
	//if (out_en101 == 1'd1) $fwrite(my_output, "%d\n", io_out101);
	//if (out_en102 == 1'd1) $fwrite(my_output, "%d\n", io_out102);
	//if (out_en103 == 1'd1) $fwrite(my_output, "%d\n", io_out103);
	//if (out_en104 == 1'd1) $fwrite(my_output, "%d\n", io_out104);
	//if (out_en105 == 1'd1) $fwrite(my_output, "%d\n", io_out105);
	//if (out_en106 == 1'd1) $fwrite(my_output, "%d\n", io_out106);
	//if (out_en107 == 1'd1) $fwrite(my_output, "%d\n", io_out107);
	//if (out_en108 == 1'd1) $fwrite(my_output, "%d\n", io_out108);
	//if (out_en109 == 1'd1) $fwrite(my_output, "%d\n", io_out109);
	//if (out_en110 == 1'd1) $fwrite(my_output, "%d\n", io_out110);
	//if (out_en111 == 1'd1) $fwrite(my_output, "%d\n", io_out111);
	//if (out_en112 == 1'd1) $fwrite(my_output, "%d\n", io_out112);
	//if (out_en113 == 1'd1) $fwrite(my_output, "%d\n", io_out113);
	//if (out_en114 == 1'd1) $fwrite(my_output, "%d\n", io_out114);
	//if (out_en115 == 1'd1) $fwrite(my_output, "%d\n", io_out115);
	//if (out_en116 == 1'd1) $fwrite(my_output, "%d\n", io_out116);
	//if (out_en117 == 1'd1) $fwrite(my_output, "%d\n", io_out117);
	//if (out_en118 == 1'd1) $fwrite(my_output, "%d\n", io_out118);
	//if (out_en119 == 1'd1) $fwrite(my_output, "%d\n", io_out119);
	//if (out_en120 == 1'd1) $fwrite(my_output, "%d\n", io_out120);
	//if (out_en121 == 1'd1) $fwrite(my_output, "%d\n", io_out121);
	//if (out_en122 == 1'd1) $fwrite(my_output, "%d\n", io_out122);
	//if (out_en123 == 1'd1) $fwrite(my_output, "%d\n", io_out123);
	//if (out_en124 == 1'd1) $fwrite(my_output, "%d\n", io_out124);
	//if (out_en125 == 1'd1) $fwrite(my_output, "%d\n", io_out125);
	//if (out_en126 == 1'd1) $fwrite(my_output, "%d\n", io_out126);
	//if (out_en127 == 1'd1) $fwrite(my_output, "%d\n", io_out127);
	//if (out_en128 == 1'd1) $fwrite(my_output, "%d\n", io_out128);
	//if (out_en129 == 1'd1) $fwrite(my_output, "%d\n", io_out129);
	//if (out_en130 == 1'd1) $fwrite(my_output, "%d\n", io_out130);
	//if (out_en131 == 1'd1) $fwrite(my_output, "%d\n", io_out131);
	//if (out_en132 == 1'd1) $fwrite(my_output, "%d\n", io_out132);
	//if (out_en133 == 1'd1) $fwrite(my_output, "%d\n", io_out133);
	//if (out_en134 == 1'd1) $fwrite(my_output, "%d\n", io_out134);
	//if (out_en135 == 1'd1) $fwrite(my_output, "%d\n", io_out135);
	//if (out_en136 == 1'd1) $fwrite(my_output, "%d\n", io_out136);
	//if (out_en137 == 1'd1) $fwrite(my_output, "%d\n", io_out137);
	//if (out_en138 == 1'd1) $fwrite(my_output, "%d\n", io_out138);
	//if (out_en139 == 1'd1) $fwrite(my_output, "%d\n", io_out139);
end



multicore multicore(clk, in, io_out0, io_out1,// io_out2, io_out3, io_out4, io_out5, io_out6, io_out7, io_out8, io_out9, io_out10, io_out11, io_out12, io_out13, io_out14, io_out15, io_out16, io_out17, io_out18, io_out19, io_out20, io_out21, io_out22, io_out23, io_out24, io_out25, io_out26, io_out27, io_out28, io_out29, io_out30, io_out31, io_out32, io_out33, io_out34, io_out35, io_out36, io_out37, io_out38, io_out39, io_out40, io_out41, io_out42, io_out43, io_out44, io_out45, io_out46, io_out47, io_out48, io_out49, io_out50, io_out51, io_out52, io_out53, io_out54, io_out55, io_out56, io_out57, io_out58, io_out59, io_out60, io_out61, io_out62, io_out63, io_out64, io_out65, io_out66, io_out67, io_out68, io_out69, io_out70, io_out71, io_out72, io_out73, io_out74, io_out75, io_out76, io_out77, io_out78, io_out79, io_out80, io_out81, io_out82, io_out83, io_out84, io_out85, io_out86, io_out87, io_out88, io_out89, io_out90, io_out91, io_out92, io_out93, io_out94, io_out95, io_out96, io_out97, io_out98, io_out99, io_out100, io_out101, io_out102, io_out103, io_out104, io_out105, io_out106, io_out107, io_out108, io_out109, io_out110, io_out111, io_out112, io_out113, io_out114, io_out115, io_out116, io_out117, io_out118, io_out119, io_out120, io_out121, io_out122, io_out123, io_out124, io_out125, io_out126, io_out127, io_out128, io_out129, io_out130, io_out131, io_out132, io_out133, io_out134, io_out135, io_out136, io_out137, io_out138, io_out139, 
req_in0, req_in1,// req_in2, req_in3, req_in4, req_in5, req_in6, req_in7, req_in8, req_in9, req_in10, req_in11, req_in12, req_in13, req_in14, req_in15, req_in16, req_in17, req_in18, req_in19, req_in20, req_in21, req_in22, req_in23, req_in24, req_in25, req_in26, req_in27, req_in28, req_in29, req_in30, req_in31, req_in32, req_in33, req_in34, req_in35, req_in36, req_in37, req_in38, req_in39, req_in40, req_in41, req_in42, req_in43, req_in44, req_in45, req_in46, req_in47, req_in48, req_in49, req_in50, req_in51, req_in52, req_in53, req_in54, req_in55, req_in56, req_in57, req_in58, req_in59, req_in60, req_in61, req_in62, req_in63, req_in64, req_in65, req_in66, req_in67, req_in68, req_in69, req_in70, req_in71, req_in72, req_in73, req_in74, req_in75, req_in76, req_in77, req_in78, req_in79, req_in80, req_in81, req_in82, req_in83, req_in84, req_in85, req_in86, req_in87, req_in88, req_in89, req_in90, req_in91, req_in92, req_in93, req_in94, req_in95, req_in96, req_in97, req_in98, req_in99, req_in100, req_in101, req_in102, req_in103, req_in104, req_in105, req_in106, req_in107, req_in108, req_in109, req_in110, req_in111, req_in112, req_in113, req_in114, req_in115, req_in116, req_in117, req_in118, req_in119, req_in120, req_in121, req_in122, req_in123, req_in124, req_in125, req_in126, req_in127, req_in128, req_in129, req_in130, req_in131, req_in132, req_in133, req_in134, req_in135, req_in136, req_in137, req_in138, req_in139,
out_en0, out_en1);//, out_en2, out_en3, out_en4, out_en5, out_en6, out_en7, out_en8, out_en9, out_en10, out_en11, out_en12, out_en13, out_en14, out_en15, out_en16, out_en17, out_en18, out_en19, out_en20, out_en21, out_en22, out_en23, out_en24, out_en25, out_en26, out_en27, out_en28, out_en29, out_en30, out_en31, out_en32, out_en33, out_en34, out_en35, out_en36, out_en37, out_en38, out_en39, out_en40, out_en41, out_en42, out_en43, out_en44, out_en45, out_en46, out_en47, out_en48, out_en49, out_en50, out_en51, out_en52, out_en53, out_en54, out_en55, out_en56, out_en57, out_en58, out_en59, out_en60, out_en61, out_en62, out_en63, out_en64, out_en65, out_en66, out_en67, out_en68, out_en69, out_en70, out_en71, out_en72, out_en73, out_en74, out_en75, out_en76, out_en77, out_en78, out_en79, out_en80, out_en81, out_en82, out_en83, out_en84, out_en85, out_en86, out_en87, out_en88, out_en89, out_en90, out_en91, out_en92, out_en93, out_en94, out_en95, out_en96, out_en97, out_en98, out_en99, out_en100, out_en101, out_en102, out_en103, out_en104, out_en105, out_en106, out_en107, out_en108, out_en109, out_en110, out_en111, out_en112, out_en113, out_en114, out_en115, out_en116, out_en117, out_en118, out_en119, out_en120, out_en121, out_en122, out_en123, out_en124, out_en125, out_en126, out_en127, out_en128, out_en129, out_en130, out_en131, out_en132, out_en133, out_en134, out_en135, out_en136, out_en137, out_en138, out_en139);

endmodule
